LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY display IS
PORT (  clk2 : IN STD_LOGIC;
        CQIN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        CQHigh:in STD_LOGIC_VECTOR(15 downto 0);
        SG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
        BT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) );
END;
ARCHITECTURE one OF display IS
SIGNAL CNT8 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL A:STD_LOGIC_VECTOR(3 downto 0);
SIGNAL B:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL COUNT:STD_LOGIC_VECTOR(9 DOWNTO 0):="0000000000";
SIGNAL CLK3:STD_LOGIC:='0';
BEGIN

P0:PROCESS(CLK2)
BEGIN

    IF CLK2 ='1' AND CLK2'EVENT
        THEN
        COUNT<=COUNT+'1';
        IF COUNT="1111111111"
        THEN CLK3<=NOT CLK3;
        COUNT<="0000000000";
        END IF;
     END IF;



END PROCESS P0;

P1: PROCESS( CNT8 )
BEGIN
CASE CNT8 IS
WHEN "000" => BT <= "11111110" ; A <= CQIN(3 DOWNTO 0) ;
WHEN "001" => BT <= "11111101" ; A <=CQIN(7 DOWNTO 4) ;
WHEN "010" => BT <= "11111011" ; A <= CQIN(11 DOWNTO 8) ;
WHEN "011" => BT <= "11110111" ; A <= CQIN(15 DOWNTO 12) ;
WHEN "100" => BT <= "11101111" ; A <= CQHigh(3 DOWNTO 0) ;
WHEN "101" => BT <= "11011111" ; A <= CQHigh(7 DOWNTO 4) ;
WHEN "110" => BT <= "10111111" ; A <= CQHigh(11 DOWNTO 8) ;
WHEN "111" => BT <= "01111111" ; A <= CQHigh(15 DOWNTO 12) ;
WHEN OTHERS => NULL ;
END CASE ;
END PROCESS P1;

P2: PROCESS(CLK3)
BEGIN
IF CLK3'EVENT AND CLK3 = '1' THEN CNT8 <= CNT8 + '1';
END IF;
END PROCESS P2 ;
P3: PROCESS(A) --�����·
BEGIN
CASE A IS
WHEN "0000" => SG <= "11000000"; WHEN "0001" => SG <= "11111001";
WHEN "0010" => SG <= "10100100"; WHEN "0011" => SG <= "10110000";
WHEN "0100" => SG <= "10011001"; WHEN "0101" => SG <= "10010010";
WHEN "0110" => SG <= "10000010"; WHEN "0111" => SG <= "11111000";
WHEN "1000" => SG <= "10000000"; WHEN "1001" => SG <= "10010000";
WHEN "1010" => SG <= "10001000"; WHEN "1011" => SG <= "10000011";
WHEN "1100" => SG <= "11000110"; WHEN "1101" => SG <= "10100001";
WHEN "1110" => SG <= "10000110"; WHEN "1111" => SG <= "10001110";

WHEN OTHERS => NULL ;
END CASE ;
END PROCESS P3;
END;
